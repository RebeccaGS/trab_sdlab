entity complement_2 is
    port (
        A         : in  STD_LOGIC_VECTOR(3 downto 0); -- A0 A1 A2 A3
        Z         : out STD_LOGIC_VECTOR(3 downto 0);
    );
end entity complement_2;